`define WIDTH 8
`define DEPTH 8
